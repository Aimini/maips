typedef struct {
    compare_t compare;
    logic carry,overflow;
} flag_t;