module stage_memory_test();
    

endmodule