typedef struct {
    compare_t compare;
    logic carry;
} flag_t;