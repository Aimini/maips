typedef  struct {
    logic eq,neq,gt,lt,gtu,ltu;
} compare_t;