`include "src/top.sv"

module top_test();
    logic clk,reset;

    always begin
        clk = 1; #5ns;
        clk = 0; #5ns;
    end

    top unit_top(clk,reset);

    logic[31:0] reg_v[1:0],reg_a[3:0],reg_s[7:0],reg_t[9:0];
    logic[31:0]  reg_file[31:0];
    logic write_dbg_memory;
    logic[31:0] dbg_arg[7:0];
    logic[31:0] previous_dbg_arg;

    string dbg_target = "sw_dbg";
    string target_name[] = '{dbg_target,"lui","ori"};
    string test_target = target_name[1];
    string test_file = {"asm/temp/", test_target, ".asm.hextext"};
    string regchk_file = {"asm/temp/", test_target, ".reg.hextext"};

    always_comb begin
        reg_file = unit_top.unit_core.unit_decode.unit_rf.file;
        reg_v  =  reg_file[3:2];
        reg_a  = reg_file[7:4];
        reg_s = reg_file[23:16];
        reg_t = {reg_file[25:24], reg_file[15:8]};

        write_dbg_memory =  unit_top.unit_memory.debug_we;
        dbg_arg = unit_top.unit_memory.unit_debug_ram.datas;
    end

    /* fill for sw_dbg test */
    task fill_regsiter_sw_dbg();
       unit_top.unit_core
       .unit_decode.unit_rf.file[2] = 32'hffff0000; //v0 = 0xFFFF0000
       for(int i = 0; i < 8; ++i)
            unit_top.unit_core
            .unit_decode.unit_rf.file[16 + i] =  1 << i; //s0 - s7
        unit_top.unit_core
       .unit_decode.unit_rf.file[16] = 32'hffff0000; //s0 = 0xFFFF0000
    endtask
    
    /** check reg file **/
    function automatic void check_regfile(string filename,logic[31:0]  rf[31:0],logic ignore_gp_sp);
        logic[31:0]  temp[31:0];
        $readmemh(regchk_file, temp);
            for(int i = 0; i < 32; ++i) begin
                if(ignore_gp_sp & (i == 28 | i == 29))
                    continue;
                assert (temp[i] === rf[i]) 
                else   $error("register file check failed at %0d: %8h != %8h ",i,temp[i],rf[i]);
            end
    endfunction;


    initial begin
        reset = 1;

        $readmemh(test_file, unit_top.unit_memory.unit_ins_rom.im);
        @(negedge clk) begin
            reset = 1;
        end
        
        @(negedge clk) begin
            if(test_target == dbg_target) begin
                fill_regsiter_sw_dbg();
            end

            reset = 0;
        end
    end


    always @(negedge clk) begin
        if(previous_dbg_arg !== dbg_arg[0])  begin
            case(dbg_arg[0])
                0: $finish;

                1: begin
                    assert(dbg_arg[1] !== dbg_arg[2])
                    else $error("assert equal failed : %8h != %8h",dbg_arg[1],dbg_arg[2]);
                end

                2:  begin
                    assert(dbg_arg[1] !== dbg_arg[2])
                    else $error("assert not equal failed : %8h == %8h",dbg_arg[1],dbg_arg[2]);
                end

                // check regiter file with pattern
                // 32'h0005_0000 32'h000A_0000 32'h0014_0000 32'h0028_0000
                // 32'h0050_0000 32'h00A0_0000 32'h0140_0000 32'h0280_0000 and so on
                32'h0001_0000: begin
                    if(dbg_arg[1] === 32'h0001_0000)
                        check_regfile(regchk_file,reg_file,1);
                    else
                        check_regfile(regchk_file,reg_file,0);
                end

                32'hffff_0000: begin
                    for(int i = 0; i < 8; ++i) begin
                        $display("dbg(%0d) = %8h",i,dbg_arg[i]);
                    end
                    // check dbg_arg memory 
                    if(dbg_arg[1] == 32'h0000_0020) begin
                        assert (dbg_arg[0] === 32'hffff_0000)
                        else  $error("dbg(0) != 32'hffff_0000!");
                        for(int i = 1; i < 8; ++i) begin
                            assert (dbg_arg[i] === (1 << i))
                            else  $error("sw_dbg failed: dbg(%0d) != %8h",i,dbg_arg[i]);
                        end
                    end
                end

                default:
                    $error("unsupport check!");
            endcase
        end
        previous_dbg_arg = dbg_arg[0];
    end
endmodule