typedef struct {
    compare_t compare;
    logic rt_zero;
} flag_t;